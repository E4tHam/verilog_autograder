
module or_gate (
    input a, b,
    output wire c
);

    assign c = a || b;

endmodule
